module comms (
    input clk,
    input 
