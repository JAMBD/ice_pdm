module comms_testbench;
endmodule
