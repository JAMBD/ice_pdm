module top (
        input RX,
        output TX,
);

assign TX = RX;
endmodule

